library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity prec_add is
  generic(
    B    :   integer := 16;
    L    :   integer := 4
    );
    port(
      i_theta_H : in signed(0 to B-L);
      sigma : in std_logic_vector(0 to L-1);
      o_theta_H : out signed(0 to B-L)
    );
end entity prec_add;

architecture beh of prec_add is

  type E_TABLE is array (0 to L-1) of signed(0 to B-L);
  signal e : E_TABLE:=("000000110100100011100111101111101010000101010","000000011001000101001000100000101100101101110","000001011001010111111100101000100101011101111","000010001001000110100110010110101011101110000","000000100100010001010110100010100001001011011","000001010101001000100010010001101011110111000","000000101010101010010001000100010100111101000","000000010101010101010100100010001000000011111","000000000010101010101010101001000100001111100","000000000000010101010101010101010010001001000","000000000000000010101010101010101010100100001","000000000000000000010101010101010101010101001","000000000000000000000010101010101010101010101","000000000000000000000000010101010101010101010","000000000000000000000000000010101010101010101","000000000000000000000000000000010101010101010","000000000000000000000000000000000010101010101","000000000000000000000000000000000000010101010","000000000000000000000000000000000000000010101","000000000000000000000000000000000000000000010");

  type t_array is array (0 to L) of signed(0 to B-L);
  signal theta_arr : t_array;

begin
  
  theta_arr(0)<=i_theta_H;
  o_theta_H<=theta_arr(L)-"010000000000000000000000000000000000000000000";

  gen_add: 
   for i in 0 to L-1 generate
     theta_arr(i+1)<= theta_arr(i)+e(i) when sigma(i)='1' else
                      theta_arr(i)-e(i);
   end generate gen_add;

end architecture beh;

