library IEEE;
    use IEEE.std_logic_1164.all;
    use IEEE.numeric_std.all;
    use IEEE.fixed_float_types.all;
    use IEEE.fixed_pkg.all;
    use STD.textio.all;
    use ieee.std_logic_textio.all;
    use std.env.finish;
    
entity testbench is
    end testbench;
    
    architecture tb of testbench is
    
    component basic_cordic is
    GENERIC (
        NMB_ITERATIONS  :   integer := 30;
        PRECISION_FP    :   integer := 31
    );
    
port (
        angle_i : in sfixed (1 downto - PRECISION_FP);
        start_i : in std_logic;
        clock_i : in std_logic;
        sin_o : out sfixed (1 downto - PRECISION_FP);
        cos_o : out sfixed (1 downto - PRECISION_FP);
        rdy_o : out std_logic);
    end component;
    
component clkGen is
    port (clk : out std_logic);
    end component;
    
signal sig_clk, sig_start, sig_rdy: std_logic;
    signal sin_out, cos_out : sfixed (1 downto -31);
    signal sig_in : sfixed (1 downto -31);
    

begin
       
    -- connect DUT with tb signals
    DUT:
        basic_cordic
        generic map(NMB_ITERATIONS => 30, PRECISION_FP => 31)
        port map(
        angle_i => sig_in,
        start_i => sig_start,
        clock_i => sig_clk,
        rdy_o => sig_rdy,
        sin_o => sin_out,
        cos_o => cos_out);
            
    -- clockgenerator
    mClkGen : clkGen port map(
        clk => sig_clk
    );
        
    -- apply a test angle as input
    stimuli: process
    begin
        sig_in <= to_sfixed(-0.7853981633974483, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(-0.7696902001294993, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(-0.7539822368615503, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(-0.7382742735936014, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(-0.7225663103256524, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(-0.7068583470577035, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(-0.6911503837897545, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(-0.6754424205218055, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(-0.6597344572538566, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(-0.6440264939859076, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(-0.6283185307179586, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(-0.6126105674500096, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(-0.5969026041820606, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(-0.5811946409141118, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(-0.5654866776461627, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(-0.5497787143782138, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(-0.5340707511102648, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(-0.5183627878423158, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(-0.5026548245743669, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(-0.4869468613064179, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(-0.47123889803846897, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(-0.45553093477052, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(-0.439822971502571, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(-0.42411500823462206, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(-0.40840704496667307, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(-0.3926990816987241, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(-0.37699111843077515, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(-0.36128315516282616, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(-0.3455751918948772, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(-0.32986722862692824, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(-0.31415926535897926, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(-0.2984513020910303, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(-0.28274333882308134, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(-0.26703537555513235, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(-0.25132741228718336, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(-0.23561944901923448, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(-0.2199114857512855, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(-0.2042035224833365, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(-0.18849555921538752, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(-0.17278759594743853, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(-0.15707963267948966, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(-0.14137166941154067, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(-0.12566370614359168, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(-0.10995574287564269, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(-0.0942477796076937, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(-0.07853981633974472, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(-0.06283185307179584, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(-0.04712388980384685, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(-0.031415926535897865, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(-0.015707963267948877, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(1.1102230246251565e-16, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(0.015707963267948988, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(0.031415926535897976, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(0.04712388980384696, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(0.06283185307179595, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(0.07853981633974494, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(0.09424777960769393, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(0.1099557428756428, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(0.1256637061435918, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(0.14137166941154078, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(0.15707963267948977, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(0.17278759594743875, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(0.18849555921538763, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(0.20420352248333662, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(0.2199114857512856, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(0.23561944901923448, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(0.2513274122871836, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(0.26703537555513246, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(0.28274333882308156, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(0.29845130209103043, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(0.3141592653589793, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(0.3298672286269284, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(0.3455751918948773, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(0.3612831551628264, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(0.37699111843077526, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(0.39269908169872414, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(0.40840704496667324, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(0.4241150082346221, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(0.4398229715025712, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(0.4555309347705201, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(0.47123889803846897, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(0.48694686130641807, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(0.5026548245743669, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(0.518362787842316, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(0.5340707511102649, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(0.549778714378214, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(0.5654866776461629, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(0.5811946409141118, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(0.5969026041820609, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(0.6126105674500097, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(0.6283185307179588, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(0.6440264939859077, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(0.6597344572538566, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(0.6754424205218057, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(0.6911503837897546, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(0.7068583470577037, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(0.7225663103256525, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(0.7382742735936014, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(0.7539822368615505, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
        sig_in <= to_sfixed(0.7696902001294994, 1, - 31);
        sig_start <= '1';
        wait until sig_rdy = '1';
        sig_start <= '0';
        std.textio.write(std.textio.output, to_string(cos_out) & LF);
        std.textio.write(std.textio.output, to_string(sin_out) & LF);
        wait for 20 ns;
   finish;
    end process stimuli;
end;

